//////////////////////////////////////////////////////////////////////////////////
// Exercise #7
// Student Name: Devang Sehgal
// Date: 11 June 2020
//
//  Description: In this exercise, you need to implement a times table of 0..7x0..7
//  using a memory.
//
//  inputs:
//           clk, a[2:0], b[2:0], read
//
//  outputs:
//           result[4:0]
// edit: should be result[5:0]
//////////////////////////////////////////////////////////////////////////////////

`timescale 1ns / 100ps

module multiply(
    //Todo: add ports
    input clk,
    input [2:0] a,
    input [2:0] b,
    input read,
    output [5:0] result
    );


    //Todo: define registers and wires here

    //Todo: define your logic here


endmodule
