//////////////////////////////////////////////////////////////////////////////////
// Exercise #8
// Student Name: Devang Sehgal
// Date: 11 June 2020
//
//  Description: In this exercise, you need to implement a times table of 0..7x0..7
//  using a memory and AXI-4-lite interface.
//
//  inputs:
//           clk, rst, a[2:0], b[2:0], enable
//
//  outputs:
//           result[5:0]
//////////////////////////////////////////////////////////////////////////////////

`timescale 1ns / 100ps

module multiply_2(
    //Todo: add ports
    input clk,
    input rst,
    input [2:0] a,
    input [2:0] b,
    input enable,
    output [5:0] result
    );


    //Todo: define registers and wires here




endmodule
